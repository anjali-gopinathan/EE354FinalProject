`timescale 1ns / 1ps

module block_controller(
	input clk, //this clock must be a slow enough clock to view the changing positions of the objects
	input bright,
	input rst,
	input up, input down, input left, input right,
	input [9:0] hCount, vCount,
	output reg [11:0] rgb,
	output reg [11:0] background
   );
	wire paddle_fill;

	integer block_grid_i, integer block_grid_j;
	integer i = 0;
	
	//these two values dictate the center of the block, incrementing and decrementing them leads the block to move in certain directions
	reg [9:0] xpos, ypos;
	
	parameter RED   = 12'b1111_0000_0000;
	parameter PINK  = 12'b1111_0000_1111;
	
/**	Fill grid of blocks
*/	
	// reg [60:0] blocks;
	reg [12:0] blocks [60:0];

	// each block will be 53 wide, 12 blocks wide, 0px in between each block
	// 25 pixels tall, 5 rows, 0 px in between

	for( block_grid_i = 0; block_grid_i < 5; block_grid_i++ ){		// i represents rows
		for(block_grid_j = 0; block_grid_j < 12; block_grid_j++){		
			// assign paddle_fill=vCount>=(ypos-5) && vCount<=(ypos+5) && hCount>=(xpos-25) && hCount<=(xpos+25);
			
			// currently not storing coordinates, but assigning blocks to spots. need to store these in an 
			// array later but idk how to do that yet so we're j overwriting the same variable 
			assign blocks[i] = 
				vCount >= ((block_grid_i*25) + 50) &&		// top
				vCount <= ((block_grid_i*25) + 75) &&		// bottom
				hCount >= ((block_grid_j*53) + 150) &&		// left
				hCount <= ((block_grid_j*53) + 203);		// right
			i <= i + 1;
		}
	}

	/*when outputting the rgb value in an always block like this, make sure to include the if(~bright) statement, as this ensures the monitor 
	will output some data to every pixel and not just the images you are trying to display*/
	always@ (*) begin
    	if(~bright )	//force black if not inside the display area
			rgb = 12'b0000_0000_0000;
		else if (paddle_fill) 
			rgb = RED; 
		else if (blocks)
			rgb = PINK;
		else	
			rgb=background;
	end
		//the +-5 for the positions give the dimension of the block (i.e. it will be 50x10 pixels), 50 wide, 10 tall
	assign paddle_fill=vCount>=(ypos-5) && vCount<=(ypos+5) && hCount>=(xpos-25) && hCount<=(xpos+25);
	
	always@(posedge clk, posedge rst) 
	begin
		if(rst)
		begin 
			//rough values for center of screen
			xpos<=450;
			ypos<=500;
		end
		else if (clk) begin
		
		/* Note that the top left of the screen does NOT correlate to vCount=0 and hCount=0. The display_controller.v file has the 
			synchronizing pulses for both the horizontal sync and the vertical sync begin at vcount=0 and hcount=0. Recall that after 
			the length of the pulse, there is also a short period called the back porch before the display area begins. So effectively, 
			the top left corner corresponds to (hcount,vcount)~(144,35). Which means with a 640x480 resolution, the bottom right corner 
			corresponds to ~(783,515).  
		*/
			if(right) begin
				xpos<=xpos+2; //change the amount you increment to make the speed faster 
				if(xpos==800) //these are rough values to attempt looping around, you can fine-tune them to make it more accurate- refer to the block comment above
					xpos<=800;		// if wrapping, set to 150
			end
			else if(left) begin
				xpos<=xpos-2;
				if(xpos==150)
					xpos<=150;		// if wrapping, set xpos to 800
			end
			// else if(up) begin
			// 	ypos<=ypos-2;
			// 	if(ypos==34)
			// 		ypos<=514;
			// end
			// else if(down) begin
			// 	ypos<=ypos+2;
			// 	if(ypos==514)
			// 		ypos<=34;
			// end
		end
	end
	
	//the background color reflects the most recent button press
	always@(posedge clk, posedge rst) begin
		// if(rst)
		background <= 12'b1111_1111_1111;
		// else 
		// 	if(right)
		// 		background <= 12'b1111_1111_0000;		// yellow orange ish
		// 	else if(left)
		// 		background <= 12'b0000_1111_1111;		// light blue
		// 	else if(down)
		// 		background <= 12'b0000_1111_0000;		// bright green
		// 	else if(up)
		// 		background <= 12'b0000_0000_1111;		// royal blue
	end

	
	
endmodule
